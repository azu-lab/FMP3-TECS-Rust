signature sTaskBody {
	void main(void);
};

[active, generate(RustFMP3Plugin, "TASK, lib")]
celltype tTaskRs {
	call	sTaskBody	cTaskBody;

	attr {
		[omit] PLType("ID")				id = PL_EXP("TSKID_$id$");
		PLType("itron::task::TaskRef<'static>")			task_ref = PL_EXP("unsafe{itron::task::TaskRef::from_raw_nonnull(NonZeroI32::new(TSKID_$id$).unwrap())}");
		[omit] PLType("ATR")		attribute = PL_EXP("TA_NULL");
		[omit] PLType("PRI")		priority = PL_EXP("0");
		[omit] PLType("size_t")	stackSize = PL_EXP("0");
		[omit] PLType("size_t")	systemStackSize = PL_EXP("0");
	};
};