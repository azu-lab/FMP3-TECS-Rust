/*
 *  カーネルオブジェクトの定義
 */

signature sCheck {
    uint32_t add([in] uint32_t i, [in] uint32_t j);
    void sub([in] int32_t i, [in] int32_t j, [out] int32_t* result);
    int32_t sum([in, size_is(8)] const int32_t* array);
    void copy([in, size_is(8)] const int32_t* input, [out, size_is(8)] int32_t** output);
};

[generate(RustASP3CelltypePlugin, "lib")]
celltype tRustCall{
    call sCheck cEntry;
    entry sCheck eRustCall;
    attr {
        uint32_t id = 0;
    };
};

[generate(RustASP3CelltypePlugin, "lib")]
celltype tRustEntry{
    entry sCheck eRustEntry;
    attr {
        uint32_t id = 0;
    };
};

celltype tCCall{
    call sCheck cEntry;
    entry sCheck eCEntry;
    attr {
        uint32_t id = 0;
    };
};

celltype tCEntry{
    entry sCheck eCEntry;
    attr {
        uint32_t id = 0;
    };
};


// Rust-C
cell tRustCall RustCall {
    cEntry = CEntry.eCEntry;
    id = 0;
};
cell tCEntry CEntry {
    id = 1;
};

// C-Rust
cell tCCall CCall {
    cEntry = RustEntry.eRustEntry;
    id = 0;
};
cell tRustEntry RustEntry {
    id = 1;
};

// Rust-Rust 
cell tRustCall RustCall2 {
    cEntry = RustEntry.eRustEntry;
    id = 0;
};

// C-C
cell tCCall CCall2 {
    cEntry = CEntry.eCEntry;
    id = 0;
};