/*
 *  TOPPERS/FMP Kernel
 *      Toyohashi Open Platform for Embedded Real-Time Systems/
 *      Multi-Processor
 * 
 *  Copyright (C) 2015,2016 by Ushio Laboratory
 *              Graduate School of Engineering Science, Osaka Univ., JAPAN
 *  Copyright (C) 2015-2018 by Embedded and Real-Time Systems Laboratory
 *              Graduate School of Information Science, Nagoya Univ., JAPAN
 *  Copyright (C) 2019 by TOPPERS Project
 * 
 *  上記著作権者は，以下の(1)〜(4)の条件を満たす場合に限り，本ソフトウェ
 *  ア（本ソフトウェアを改変したものを含む．以下同じ）を使用・複製・改
 *  変・再配布（以下，利用と呼ぶ）することを無償で許諾する．
 *  (1) 本ソフトウェアをソースコードの形で利用する場合には，上記の著作
 *      権表示，この利用条件および下記の無保証規定が，そのままの形でソー
 *      スコード中に含まれていること．
 *  (2) 本ソフトウェアを，ライブラリ形式など，他のソフトウェア開発に使
 *      用できる形で再配布する場合には，再配布に伴うドキュメント（利用
 *      者マニュアルなど）に，上記の著作権表示，この利用条件および下記
 *      の無保証規定を掲載すること．
 *  (3) 本ソフトウェアを，機器に組み込むなど，他のソフトウェア開発に使
 *      用できない形で再配布する場合には，次のいずれかの条件を満たすこ
 *      と．
 *    (a) 再配布に伴うドキュメント（利用者マニュアルなど）に，上記の著
 *        作権表示，この利用条件および下記の無保証規定を掲載すること．
 *    (b) 再配布の形態を，別に定める方法によって，TOPPERSプロジェクトに
 *        報告すること．
 *  (4) 本ソフトウェアの利用により直接的または間接的に生じるいかなる損
 *      害からも，上記著作権者およびTOPPERSプロジェクトを免責すること．
 *      また，本ソフトウェアのユーザまたはエンドユーザからのいかなる理
 *      由に基づく請求からも，上記著作権者およびTOPPERSプロジェクトを
 *      免責すること．
 * 
 *  本ソフトウェアは，無保証で提供されているものである．上記著作権者お
 *  よびTOPPERSプロジェクトは，本ソフトウェアに関して，特定の使用目的
 *  に対する適合性も含めて，いかなる保証も行わない．また，本ソフトウェ
 *  アの利用により直接的または間接的に生じたいかなる損害に関しても，そ
 *  の責任を負わない．
 * 
 *  $Id: kernel.cdl 285 2018-03-21 02:55:49Z ertl-hiro $
 */

/*
 *		TOPPERS/FMPカーネルオブジェクト コンポーネント記述ファイル
 */

/*
 *  カーネルオブジェクトのコンポーネント化のためのヘッダファイル
 */
import_C("tecs_kernel.h");

typedef	int_t	TaskRef;
//typedef	int_t	MutexRef;
typedef int_t ITRONResult__empty__ActivateError__;
typedef int_t ITRONResult__empty__ActivateOnError__;
typedef int_t ITRONResult__usize__CancelActivateAllError__;
typedef int_t ITRONResult__empty__SetPriorityError__;
typedef int_t Priority;
typedef int_t ITRONResult__Priority__PriorityError__;
typedef int_t ITRONResult__empty__MigrateError__;
typedef int_t Processor;
typedef int_t ITRONResult__State__StateError__;
typedef int_t ITRONResult__Info__InfoError__;
typedef int_t ITRONResult__empty__WakeError__;
typedef int_t ITRONResult__usize__CancelWakeAllError__;
typedef int_t ITRONResult__empty__ReleaseWaitError__;
typedef int_t ITRONResult__empty__SuspendError__;
typedef int_t ITRONResult__empty__ResumeError__;
typedef int_t ITRONResult__empty__RaiseTerminationError__;
typedef int_t ITRONResult__empty__TerminateError__;


/*
 *  タスク操作のシグニチャ（タスクコンテキスト用）
 */
signature sTaskRs {
	ITRONResult__empty__ActivateError__				activate(void);
	ITRONResult__empty__ActivateOnError__			migrateAndActivate([in] Processor prcid);           // FMP3
	ITRONResult__usize__CancelActivateAllError__	cancelActivate(void);
  	ITRONResult__empty__MigrateError__    			migrate([in] Processor prcid);                      // FMP3
	ITRONResult__State__StateError__				getTaskState(void);
	ITRONResult__empty__SetPriorityError__			changePriority([in] Priority priority);
	ER												changeSubPriority([in] uint_t subPriority);  // FMP3
	ITRONResult__Priority__PriorityError__			getPriority(void);
	ITRONResult__Info__InfoError__					refer(void);

	ITRONResult__empty__WakeError__					wakeup(void);
	ITRONResult__usize__CancelWakeAllError__		cancelWakeup(void);
	ITRONResult__empty__ReleaseWaitError__			releaseWait(void);
	ITRONResult__empty__SuspendError__				suspend(void);
	ITRONResult__empty__ResumeError__				resume(void);

	ITRONResult__empty__RaiseTerminationError__		raiseTerminate(void);
	ITRONResult__empty__TerminateError__			terminate(void);
};

/*
 *  タスクのセルタイプ
 *
 *  タスクはいずれかの保護ドメインに所属させなければならない．
 */
//[active, generate(FMPObjectPlugin, "TASK"), idx_is_id]
[active, generate(FMPObjectPlugin, "TASK")]
celltype tTaskRs {
	[inline] entry	sTaskRs	eTask;
	[inline] entry	siTask	eiTask;
	call	sTaskBody	cTaskBody;

	[inline] entry	siNotificationHandler	eiActivateNotificationHandler;
	[inline] entry	siNotificationHandler	eiWakeUpNotificationHandler;

	attr {
		[omit] ID				id = C_EXP("TSKID_$id$");
		TaskRef			task_ref = C_EXP("unsafe{TaskRef::from_raw_nonnull(NonZeroI32::new(TSKID_$id$).unwrap())}");
		[omit] ATR		attribute = C_EXP("TA_NULL");
		[omit] PRI		priority;
		[omit] size_t	stackSize;
		[omit] size_t	systemStackSize = 0;
						/* 0を，未定義を示す値として使っている */
	};

	FACTORY {
		write("tecsgen.cfg", "#include \"$ct$_tecsgen.h\"");
		write("$ct$_factory.h", "#include \"kernel_cfg.h\"");
	};
};

typedef int_t SemaphoreRef;
typedef int_t ITRONResult__empty__SignalError__;
typedef int_t ITRONResult__empty__WaitError__;
typedef int_t ITRONResult__empty__PollError__;
typedef int_t ITRONResult__empty__WaitTimeoutError__;
typedef int_t Timeout;
typedef int_t ITRONResult__empty__InitializeError__;

/*
 *  セマフォ操作のシグニチャ（タスクコンテキスト用）
 */
signature sSemaphoreRs {
	ITRONResult__empty__SignalError__			signal(void);
	ITRONResult__empty__WaitError__				wait(void);
	ITRONResult__empty__PollError__				waitPolling(void);
	ITRONResult__empty__WaitTimeoutError__		waitTimeout([in] Timeout timeout);
	ITRONResult__empty__InitializeError__		initialize(void);
	ITRONResult__Info__InfoError__				refer(void);
};

/*
 *  セマフォのセルタイプ
 */
[generate(FMPObjectPlugin, "SEMAPHORE")]
celltype tSemaphoreRs {
	[inline] entry	sSemaphoreRs	eSemaphore;
	[inline] entry	siSemaphore	eiSemaphore;

	[inline] entry	siNotificationHandler	eiNotificationHandler;

	attr {
		[omit]ID				id = C_EXP("SEMID_$id$");
		SemaphoreRef	semaphore_ref = C_EXP("unsafe{SemaphoreRef::from_raw_nonnull(NonZeroI32::new(SEMID_$id$).unwrap())}");
		[omit] ATR		attribute = C_EXP("TA_NULL");
		[omit] uint_t	initialCount;
		[omit] uint_t	maxCount = 1;
	};

	FACTORY {
		write("$ct$_factory.h", "#include \"kernel_cfg.h\"");
	};
};

typedef int_t DataqueueRef;
typedef int_t ITRONResult__empty__SendError__;
typedef uint_t DataElement;
typedef int_t ITRONResult__empty__TrySendError__;
typedef int_t ITRONResult__empty__SendTimeoutError__;
typedef int_t ITRONResult__empty__SendForcedError__;
typedef int_t ITRONResult__DataElement__RecvError__;
typedef int_t ITRONResult__DataElement__TryRecvError__;
typedef int_t ITRONResult__DataElement__RecvTimeoutError__;

/*
 *  データキュー操作のシグニチャ（タスクコンテキスト用）
 */
signature sDataqueueRs {
	ITRONResult__empty__SendError__ 					send([in] DataElement data);
	ITRONResult__empty__TrySendError__ 					sendPolling([in] DataElement data);
	ITRONResult__empty__SendTimeoutError__ 				sendTimeout([in] DataElement data, [in] Timeout timeout);
	ITRONResult__empty__SendForcedError__ 				sendForce([in] DataElement data);
	ITRONResult__DataElement__RecvError__ 				receive(void);
	ITRONResult__DataElement__TryRecvError__ 			receivePolling(void);
	ITRONResult__DataElement__RecvTimeoutError__ 		receiveTimeout([in] Timeout timeout);
	ITRONResult__empty__InitializeError__ 				initialize(void);
	ITRONResult__Info__InfoError__						refer(void);
};

/*
 *  データキュー操作のシグニチャ（非タスクコンテキスト用）
 */
[context("non-task")]
signature siDataqueueRs {
	ITRONResult__empty__TrySendError__ 			sendPolling([in] DataElement data);
	ITRONResult__empty__SendForcedError__ 		sendForce([in] DataElement data);
};

/*
 *  データキューのセルタイプ
 */
[generate(FMPObjectPlugin, "DATAQUEUE")]
celltype tDataqueueRs {
	[inline] entry	sDataqueueRs	eDataqueue;
	[inline] entry	siDataqueueRs	eiDataqueue;

	[inline] entry	siNotificationHandler	eiNotificationHandler;

	attr {
		[omit] ID				id = C_EXP("DTQID_$id$");
		DataqueueRef	semaphore_ref = C_EXP("unsafe{DataqueueRef::from_raw_nonnull(NonZeroI32::new(SEMID_$id$).unwrap())}");
		[omit] ATR		attribute = C_EXP("TA_NULL");
		[omit] uint_t	dataCount = 1;
		[omit] void		*dataqueueManagementBuffer = C_EXP("NULL");
	};

	FACTORY {
		write("$ct$_factory.h", "#include \"kernel_cfg.h\"");
	};
};


// TODO: 割込みは itron_rs で実装されていないため、暫定的な実装を行う

typedef int_t ITRONResult__empty__ER__;
typedef int_t ITRONResult__bool__ER__;

/*
 *  割込み要求ライン操作のシグニチャ（タスクコンテキスト用）
 */
signature sInterruptRequestRs {
	ITRONResult__empty__ER__		disable(void);
	ITRONResult__empty__ER__		enable(void);
	ITRONResult__empty__ER__		clear(void);
	ITRONResult__empty__ER__		raise(void);
	ITRONResult__bool__ER__			probe(void);
};

/*
 *  割込み要求ラインのセルタイプ
 *
 *  割込み要求ラインはカーネルドメインに所属させなければならない．
 */
[active, generate(FMPHandlerPlugin, "INT_REQUEST")]
celltype tInterruptRequestRs {
	[inline] entry	sInterruptRequestRs	eInterruptRequest;

	attr {
		INTNO			interruptNumber;
		[omit] ATR		attribute = C_EXP("TA_NULL");
		[omit] PRI		interruptPriority;
	};

	/* 警告メッセージを抑止するための記述 */
	factory {
		write("tecsgen.cfg", "");
	};
};

/*
 *  割込みサービスルーチンのセルタイプ
 *
 */
[active, generate(FMPHandlerPlugin, "INT_SERVICE_ROUTINE")]
celltype tIsrRs {
	call	siHandlerBody	ciISRBody;

	attr {
		ID				id = C_EXP("ISRID_$id$");
		[omit] ATR		attribute = C_EXP("TA_NULL");
		[omit] INTNO	interruptNumber;
		[omit] PRI		isrPriority = 1;
	};

	FACTORY {
		write("tecsgen.cfg", "#include \"$ct$_tecsgen.h\"");
		write("$ct$_factory.h", "#include \"kernel_cfg.h\"");
	};
};